
module filter_buffer_mask_no_temp(
    );


endmodule
